library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use work.simulation_pkg.all;

package user_driver_pkg is





end user_driver_pkg;

package body user_driver_pkg is



 

end user_driver_pkg;
